`include "define.vh"

module alu (
    input wire interrupt_signal
)


endmodule
