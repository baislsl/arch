`include "define.vh"


/**
 * Data Path for MIPS 5-stage pipelined CPU.
 * Author: Zhao, Hongyu  <power_zhy@foxmail.com>
 */
module datapath (
	input wire clk,  // main clock
	// debug
	`ifdef DEBUG
	input wire [5:0] debug_addr,  // debug address
	output wire [31:0] debug_data,  // debug data
	`endif
	// control signals
    output reg mem_ren_mem,
	output reg [31:0] inst_data_id,  // instruction
	output reg [4:0] regw_addr_exe,  // register write address from EXE stage
	output reg wb_wen_exe,  // register write enable signal feedback from EXE stage
	output reg [4:0] regw_addr_mem,  // register write address from MEM stage
	output reg wb_wen_mem,  // register write enable signal feedback from MEM stage
	input wire [2:0] pc_src_ctrl,  // how would PC change to next
	input wire imm_ext_ctrl,  // whether using sign extended to immediate data
	input wire [1:0] exe_a_src_ctrl,  // data source of operand A for ALU
	input wire [1:0] exe_b_src_ctrl,  // data source of operand B for ALU
    input wire [1:0] fwd_a_ctrl,
    input wire [1:0] fwd_b_ctrl,
	input wire [3:0] exe_alu_oper_ctrl,  // ALU operation type
	input wire mem_ren_ctrl,  // memory read enable signal
	input wire mem_wen_ctrl,  // memory write enable signal
	input wire [1:0] wb_addr_src_ctrl,  // address source to write data back to registers
	input wire wb_data_src_ctrl,  // data source of data being written back to registers
	input wire wb_wen_ctrl,  // register write enable signal
	// IF signals
	input wire if_rst,  // stage reset signal
	input wire if_en,  // stage enable signal
	output reg if_valid,  // working flag
	output reg inst_ren,  // instruction read enable signal
	output reg [31:0] inst_addr,  // address of instruction needed
	input wire [31:0] inst_data,  // instruction fetched
	// ID signals
	input wire id_rst,
	input wire id_en,
	output reg id_valid,
	// EXE signals
	input wire exe_rst,
	input wire exe_en,
	output reg exe_valid,
	// MEM signals
	input wire mem_rst,
	input wire mem_en,
	output reg mem_valid,
	output wire mem_ren,  // memory read enable signal
	output wire mem_wen,  // memory write enable signal
	output wire [31:0] mem_addr,  // address of memory
	output wire [31:0] mem_dout,  // data writing to memory
	input wire [31:0] mem_din,  // data read from memory
	// WB signals
	input wire wb_rst,
	input wire wb_en,
	output reg wb_valid,
    output reg wb_wen_wb,
    output reg [4:0] regw_addr_wb,
   //rs and rd address
    output reg [4:0] addr_rs_id,// can be deleted
    output reg [4:0] addr_rs_exe,
    output reg [4:0] addr_rs_mem,
    output reg [4:0] addr_rt_id, //can be deleted
    output reg [4:0] addr_rt_exe,
    output reg [4:0] addr_rt_mem,
	 output reg [31:0] fwd_a_data,
	 output reg [31:0] fwd_b_data,
     output reg [31:0] fwd_a_data_exe,
     output reg [31:0] fwd_b_data_exe,

     output wire a_b_equal,
     input wire fwd_m,

     input wire alu_sign,

	 // interrupt
	output wire [4:0] addr_r,
	input wire [31:0] data_r,
	output wire [4:0] addr_w,
	output wire [31:0] data_w,
	output wire ir_en,
	output wire [31:0] ret_addr,
	input wire jump_en, // epc_ctrl
	input wire [31:0] jump_addr //epc
	);

	`include "mips_define.vh"

	// control signals
	reg [1:0] exe_a_src_exe, exe_b_src_exe;
	reg [3:0] exe_alu_oper_exe;
	reg mem_ren_exe;
	reg mem_wen_exe, mem_wen_mem;
	reg wb_data_src_exe, wb_data_src_mem, wb_data_src_wb;

	// IF signals
	wire [31:0] inst_addr_next;

	// ID signals
	reg [31:0] inst_addr_id;
	reg [31:0] inst_addr_next_id;
	reg [4:0] regw_addr_id;
	wire [4:0] addr_rs, addr_rt, addr_rd;
	wire [31:0] data_rs, data_rt, data_imm;

	// EXE signals
	reg [31:0] inst_addr_exe;
	reg [31:0] inst_addr_next_exe;
	reg [31:0] inst_data_exe;
	reg [31:0] data_rs_exe, data_rt_exe, data_imm_exe;
	reg [31:0] opa_exe, opb_exe;
	wire [31:0] alu_out_exe;
    reg fwd_m_exe;
	reg alu_sign_exe;
	reg [31:0] cp0_data_r_exe;

	// MEM signals
	reg [31:0] inst_addr_mem;
	reg [31:0] inst_addr_next_mem;
	reg [31:0] inst_data_mem;
	reg [31:0] data_rs_mem;	// ? [4:0] -> [31:0]
	reg [31:0] data_rt_mem;
	reg [31:0] alu_out_mem;
	reg rs_rt_equal_mem;
    reg fwd_m_mem;

	// WB signals
	reg [31:0] alu_out_wb;
	reg [31:0] mem_din_wb;
	reg [31:0] regw_data_wb;

	// debug
	`ifdef DEBUG
	wire [31:0] debug_data_reg;
	reg [31:0] debug_data_signal;

	always @(posedge clk) begin
		case (debug_addr[4:0])
			0: debug_data_signal <= inst_addr;
			1: debug_data_signal <= inst_data;
			2: debug_data_signal <= inst_addr_id;
			3: debug_data_signal <= inst_data_id;
			4: debug_data_signal <= inst_addr_exe;
			5: debug_data_signal <= inst_data_exe;
			6: debug_data_signal <= inst_addr_mem;
			7: debug_data_signal <= inst_data_mem;
			8: debug_data_signal <= {27'b0, addr_rs};
			9: debug_data_signal <= data_rs;
			10: debug_data_signal <= {27'b0, addr_rt};
			11: debug_data_signal <= data_rt;
			12: debug_data_signal <= data_imm;
			13: debug_data_signal <= opa_exe;
			14: debug_data_signal <= opb_exe;
			15: debug_data_signal <= alu_out_exe;
			16: debug_data_signal <= 0;
			17: debug_data_signal <= 0;
			18: debug_data_signal <= {19'b0, inst_ren, 7'b0, mem_ren, 3'b0, mem_wen};
			19: debug_data_signal <= mem_addr;
			20: debug_data_signal <= mem_din;
			21: debug_data_signal <= mem_dout;
			22: debug_data_signal <= {27'b0, regw_addr_wb};
			23: debug_data_signal <= regw_data_wb;
			default: debug_data_signal <= 32'hFFFF_FFFF;
		endcase
	end

	assign
		debug_data = debug_addr[5] ? debug_data_signal : debug_data_reg;
	`endif

	// IF stage
	assign
		inst_addr_next = inst_addr + 4;

	always @(*) begin
		if_valid = ~if_rst & if_en;
		inst_ren = ~if_rst;
	end

    //next PC
	always @(posedge clk) begin
		if (if_rst) begin
			inst_addr <= 0;	
		end
		else if (if_en) begin
			if(jump_en) begin
				inst_addr <= jump_addr;
			end else begin 
				case (pc_src_ctrl)
					PC_NEXT: inst_addr<=inst_addr_next;
					PC_FWD_DATA: inst_addr<=fwd_a_data;
					PC_JUMP: inst_addr<={inst_addr_id[31:28],inst_data_id[25:0], 2'b0};
					PC_BRANCH: inst_addr<=inst_addr_next_id+(data_imm<<2);
				endcase
			end 
			// if (is_branch_mem)//TODO pc select
			// 	inst_addr <= branch_target_mem;
			// else
			// 	inst_addr <= inst_addr_next;
		end
	end

	// ID stage
	always @(posedge clk) begin
		if (id_rst) begin
			id_valid <= 0;
			inst_addr_id <= 0;
			inst_data_id <= 0;
			inst_addr_next_id <= 0;
            // addr_rs_id<=0;
            // addr_rt_id<=0;
		end
		else if (id_en) begin
			id_valid <= if_valid;
			inst_addr_id <= inst_addr;
			inst_data_id <= inst_data;
			inst_addr_next_id <= inst_addr_next;
            // addr_rs_id<=addr_rs;
            // addr_rt_id<=addr_rt;
		end
	end

	assign
		addr_rs = inst_data_id[25:21],
		addr_rt = inst_data_id[20:16],
		addr_rd = inst_data_id[15:11],
		data_imm = imm_ext_ctrl ? {{16{inst_data_id[15]}}, inst_data_id[15:0]} : {16'b0, inst_data_id[15:0]};

	always @(*) begin
		regw_addr_id = inst_data_id[15:11];
		case (wb_addr_src_ctrl)
			WB_ADDR_RD: regw_addr_id = addr_rd;
			WB_ADDR_RT: regw_addr_id = addr_rt;
			WB_ADDR_LINK: regw_addr_id = GPR_RA;
		endcase
	end

	regfile REGFILE (
		.clk(clk),
		`ifdef DEBUG
		.debug_addr(debug_addr[4:0]),
		.debug_data(debug_data_reg),
		`endif
		.addr_a(addr_rs),
		.data_a(data_rs),
		.addr_b(addr_rt),
		.data_b(data_rt),
		.en_w(wb_wen_wb),
		.addr_w(regw_addr_wb),
		.data_w(regw_data_wb)
		);

	// EXE stage
	always @(posedge clk) begin
		if (exe_rst) begin
			exe_valid <= 0;
			inst_addr_exe <= 0;
			inst_data_exe <= 0;
			inst_addr_next_exe <= 0;
			regw_addr_exe <= 0;
			exe_a_src_exe <= 0;
			exe_b_src_exe <= 0;
			data_rs_exe <= 0;
			data_rt_exe <= 0;
			data_imm_exe <= 0;
			exe_alu_oper_exe <= 0;
			mem_ren_exe <= 0;
			mem_wen_exe <= 0;
			wb_data_src_exe <= 0;
			wb_wen_exe <= 0;
            addr_rs_exe<=0;
            addr_rt_exe<=0;
            fwd_a_data_exe<=0;
            fwd_b_data_exe<=0;
			alu_sign_exe<=0;
			cp0_data_r_exe<=0;
		end
		else if (exe_en) begin
			exe_valid <= id_valid;
			inst_addr_exe <= inst_addr_id;
			inst_data_exe <= inst_data_id;
			inst_addr_next_exe <= inst_addr_next_id;
			regw_addr_exe <= regw_addr_id;
			exe_a_src_exe <= exe_a_src_ctrl;
			exe_b_src_exe <= exe_b_src_ctrl;
			data_rs_exe <= data_rs;
			data_rt_exe <= data_rt;
			data_imm_exe <= data_imm;
			exe_alu_oper_exe <= exe_alu_oper_ctrl;
			mem_ren_exe <= mem_ren_ctrl;
			mem_wen_exe <= mem_wen_ctrl;
			wb_data_src_exe <= wb_data_src_ctrl;
			wb_wen_exe <= wb_wen_ctrl;
            addr_rs_exe<=addr_rs;
            addr_rt_exe<=addr_rt;
            fwd_a_data_exe<=fwd_a_data;
            fwd_b_data_exe<=fwd_b_data;
            fwd_m_exe<=fwd_m;
			alu_sign_exe<=alu_sign;
			cp0_data_r_exe<=data_r;
		end
	end

	assign
		a_b_equal = (fwd_a_data == fwd_b_data);

	assign
		// MTC0
		data_w = fwd_b_data,
		addr_w = inst_data_id[15:11],

		// MFC0
		addr_r = inst_data_id[15:11],

		ir_en = 1,
		ret_addr = pc_src_ctrl ? inst_addr_id : inst_addr;

	always @(*) begin
		// id state
        case (fwd_a_ctrl)
            2'b00: fwd_a_data=data_rs;
            2'b01:fwd_a_data=alu_out_exe;
            2'b10:fwd_a_data=alu_out_mem;
            2'b11:fwd_a_data=mem_din;
        endcase
        case (fwd_b_ctrl)
            2'b00:fwd_b_data=data_rt;
            2'b01:fwd_b_data=alu_out_exe;
            2'b10:fwd_b_data=alu_out_mem;
            2'b11:fwd_b_data=mem_din;
        endcase

		// exe state
		case (exe_a_src_exe)
			EXE_A_FWD_DATA: opa_exe = fwd_a_data_exe;
			EXE_A_LINK: opa_exe = inst_addr_next_exe;	// JAL
			EXE_A_SHIFT: opa_exe = {27'b0,inst_data_exe[10:6]};
			EXE_A_INT: opa_exe = cp0_data_r_exe;
		endcase
		case (exe_b_src_exe)
			EXE_B_FWD_DATA: opb_exe = fwd_b_data_exe;
            EXE_B_FOUR: opb_exe = 4;
			EXE_B_IMM: opb_exe = data_imm_exe;
			EXE_B_INT: opb_exe = 0;
		endcase
	end

	alu ALU (
		.a(opa_exe),
		.b(opb_exe),
		.oper(exe_alu_oper_exe),
		.result(alu_out_exe),
        .sign(alu_sign_exe)
		);

	// MEM stage
	always @(posedge clk) begin
		if (mem_rst) begin
			mem_valid <= 0;
			inst_addr_mem <= 0;
			inst_data_mem <= 0;
			inst_addr_next_mem <= 0;
			regw_addr_mem <= 0;
			data_rs_mem <= 0;
			data_rt_mem <= 0;
			alu_out_mem <= 0;
			mem_ren_mem <= 0;
			mem_wen_mem <= 0;
			wb_data_src_mem <= 0;
			wb_wen_mem <= 0;
			rs_rt_equal_mem <= 0;
            addr_rs_mem<=0;
            addr_rt_mem<=0;
            fwd_m_mem<=0;
		end
		else if (mem_en) begin
			mem_valid <= exe_valid;
			inst_addr_mem <= inst_addr_exe;
			inst_data_mem <= inst_data_exe;
			inst_addr_next_mem <= inst_addr_next_exe;
			regw_addr_mem <= regw_addr_exe;
			//data_rs_mem <= data_rs_exe;
			data_rs_mem <= fwd_a_data_exe;
			// data_rt_mem <= data_rt_exe;
			data_rt_mem <= fwd_b_data_exe;
			alu_out_mem <= alu_out_exe;
			mem_ren_mem <= mem_ren_exe;
			mem_wen_mem <= mem_wen_exe;
			wb_data_src_mem <= wb_data_src_exe;
			wb_wen_mem <= wb_wen_exe;
            addr_rs_mem<=addr_rs_exe;
            addr_rt_mem<=addr_rt_exe;
            fwd_m_mem<=fwd_m_exe;
		end
	end

    //TODO branch_target_mem
	// always @(*) begin
	// 	case (pc_src_mem)
	// 		PC_JUMP: branch_target_mem <= {inst_addr_mem[31:28],inst_data_mem[25:0], 2'b0};
	// 		PC_JR: branch_target_mem <= data_rs_mem;
	// 		PC_BEQ: branch_target_mem <= rs_rt_equal_mem ? alu_out_mem : inst_addr_next_mem;
	// 		PC_BNE: branch_target_mem <= rs_rt_equal_mem ? inst_addr_next_mem : alu_out_mem;
	// 		default: branch_target_mem <= inst_addr_next_mem;  // will never be used
	// 	endcase
	// end

	assign
		mem_ren = mem_ren_mem,
		mem_wen = mem_wen_mem,
		mem_addr = alu_out_mem,
		mem_dout = fwd_m_mem ? regw_data_wb : data_rt_mem;

	// WB stage
	always @(posedge clk) begin
		if (wb_rst) begin
			wb_valid <= 0;
			wb_wen_wb <= 0;
			wb_data_src_wb <= 0;
			regw_addr_wb <= 0;
			alu_out_wb <= 0;
			mem_din_wb <= 0;
		end
		else if (wb_en) begin
			wb_valid <= mem_valid;
			wb_wen_wb <= wb_wen_mem;
			wb_data_src_wb <= wb_data_src_mem;
			regw_addr_wb <= regw_addr_mem;
			alu_out_wb <= alu_out_mem;
			mem_din_wb <= mem_din;
		end
	end

	always @(*) begin
		regw_data_wb = alu_out_wb;
		case (wb_data_src_wb)
			WB_DATA_ALU: regw_data_wb = alu_out_wb;
			WB_DATA_MEM: regw_data_wb = mem_din_wb;
		endcase
	end

endmodule
